module LMG (clk, 
);

input clk;







endmodule