module columnUnit (clk, bstate, ...
);

input clk;
input [?:0] bstate; // board state


endmodule