module RookMapROM(
	output reg [383:0] dataOut
);


reg signed [5:0] mem[63:0];

always@(*) begin
	dataOut[5:0] = mem[0];
	dataOut[11:6] = mem[1];
	dataOut[17:12] = mem[2];
	dataOut[23:18] = mem[3];
	dataOut[29:24] = mem[4];
	dataOut[35:30] = mem[5];
	dataOut[41:36] = mem[6];
	dataOut[47:42] = mem[7];
	dataOut[53:48] = mem[8];
	dataOut[59:54] = mem[9];
	dataOut[65:60] = mem[10];
	dataOut[71:66] = mem[11];
	dataOut[77:72] = mem[12];
	dataOut[83:78] = mem[13];
	dataOut[89:84] = mem[14];
	dataOut[95:90] = mem[15];
	dataOut[101:96] = mem[16];
	dataOut[107:102] = mem[17];
	dataOut[113:108] = mem[18];
	dataOut[119:114] = mem[19];
	dataOut[125:120] = mem[20];
	dataOut[131:126] = mem[21];
	dataOut[137:132] = mem[22];
	dataOut[143:138] = mem[23];
	dataOut[149:144] = mem[24];
	dataOut[155:150] = mem[25];
	dataOut[161:156] = mem[26];
	dataOut[167:162] = mem[27];
	dataOut[173:168] = mem[28];
	dataOut[179:174] = mem[29];
	dataOut[185:180] = mem[30];
	dataOut[191:186] = mem[31];
	dataOut[197:192] = mem[32];
	dataOut[203:198] = mem[33];
	dataOut[209:204] = mem[34];
	dataOut[215:210] = mem[35];
	dataOut[221:216] = mem[36];
	dataOut[227:222] = mem[37];
	dataOut[233:228] = mem[38];
	dataOut[239:234] = mem[39];
	dataOut[245:240] = mem[40];
	dataOut[251:246] = mem[41];
	dataOut[257:252] = mem[42];
	dataOut[263:258] = mem[43];
	dataOut[269:264] = mem[44];
	dataOut[275:270] = mem[45];
	dataOut[281:276] = mem[46];
	dataOut[287:282] = mem[47];
	dataOut[293:288] = mem[48];
	dataOut[299:294] = mem[49];
	dataOut[305:300] = mem[50];
	dataOut[311:306] = mem[51];
	dataOut[317:312] = mem[52];
	dataOut[323:318] = mem[53];
	dataOut[329:324] = mem[54];
	dataOut[335:330] = mem[55];
	dataOut[341:336] = mem[56];
	dataOut[347:342] = mem[57];
	dataOut[353:348] = mem[58];
	dataOut[359:354] = mem[59];
	dataOut[365:360] = mem[60];
	dataOut[371:366] = mem[61];
	dataOut[377:372] = mem[62];
	dataOut[383:378] = mem[63];
end

initial begin
	mem[0] = 0;
	mem[1] = 0;
	mem[2] = 0;
	mem[3] = 0;
	mem[4] = 0;
	mem[5] = 0;
	mem[6] = 0;
	mem[7] = 0;
	mem[8] = 0;
	mem[9] = 0;
	mem[10] = 0;
	mem[11] = 0;
	mem[12] = 0;
	mem[13] = 0;
	mem[14] = 0;
	mem[15] = 0;
	mem[16] = 0;
	mem[17] = 0;
	mem[18] = 0;
	mem[19] = 0;
	mem[20] = 0;
	mem[21] = 0;
	mem[22] = 0;
	mem[23] = 0;
	mem[24] = 0;
	mem[25] = 0;
	mem[26] = 0;
	mem[27] = 0;
	mem[28] = 0;
	mem[29] = 0;
	mem[30] = 0;
	mem[31] = 0;
	mem[32] = 0;
	mem[33] = 0;
	mem[34] = 0;
	mem[35] = 0;
	mem[36] = 0;
	mem[37] = 0;
	mem[38] = 0;
	mem[39] = 0;
	mem[40] = 0;
	mem[41] = 0;
	mem[42] = 0;
	mem[43] = 0;
	mem[44] = 0;
	mem[45] = 0;
	mem[46] = 0;
	mem[47] = 0;
	mem[48] = 0;
	mem[49] = 0;
	mem[50] = 0;
	mem[51] = 0;
	mem[52] = 0;
	mem[53] = 0;
	mem[54] = 0;
	mem[55] = 0;
	mem[56] = 0;
	mem[57] = 0;
	mem[58] = 0;
	mem[59] = 0;
	mem[60] = 0;
	mem[61] = 0;
	mem[62] = 0;
	mem[63] = 0;
end

endmodule
